LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIVISOR IS 
PORT 
( 
CLK_IN: IN STD_LOGIC;
CLK_OUT : OUT STD_LOGIC
);
END DIVISOR;


ARCHITECTURE DIVISOR_DE_FREQ OF DIVISOR IS 
SIGNAL CONTADOR : STD_LOGIC_VECTOR (1 DOWNTO 0);
BEGIN 
PROCESS (CLK_IN)
BEGIN
IF(CLK_IN'EVENT AND CLK_IN ='1') THEN

--DISEÑO DEL CONTADOR 

   CONTADOR <= CONTADOR + "01";
	
--DISEÑO DEL COMPARADOR

   IF (CONTADOR = "11") THEN 
		CLK_OUT <= '1';
	ELSE 
		CLK_OUT <= '0';
   END IF;	
END IF;
END PROCESS;
END DIVISOR_DE_FREQ;