LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIVISOR IS 
PORT 
( 
SALIDA: BUFFER STD_LOGIC;
CLK_IN: IN STD_LOGIC
);
END DIVISOR;


ARCHITECTURE DIVISOR_DE_FREQ OF DIVISOR IS
CONSTANT TOP: STD_LOGIC_VECTOR (27 DOWNTO 0) := x"000C34F"; 
SIGNAL CONTADOR : STD_LOGIC_VECTOR (27 DOWNTO 0) := x"0000000";
SIGNAL CLK_OUT: STD_LOGIC;
BEGIN 
PROCESS (CLK_IN)
BEGIN
	IF(CLK_IN'EVENT AND CLK_IN ='1') THEN

	--DISEÑO DEL CONTADOR
	 
	  IF (CONTADOR = TOP) THEN 
	  CONTADOR <= x"0000000";
	  ELSE 
		CONTADOR <= CONTADOR + x"0000001";
	  END IF;
	  
	--DISEÑO DEL COMPARADOR

		IF (CONTADOR = TOP) THEN 
			SALIDA <= '1';
		ELSE 
			SALIDA <= '0';
		END IF;	
	END IF;
END PROCESS;


END DIVISOR_DE_FREQ;